
module TRIVIUM_CORE ( SYS_CLK, CNTRL, KEY, IV, KEY_OUT );
  input [1:0] CNTRL;
  input [79:0] KEY;
  input [79:0] IV;
  input SYS_CLK;
  output KEY_OUT;
  wire   t3, t1, t2, N301, N303, N305, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10,
         n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n750, n752, n753, n754,
         n755, n25, n110, n111, n112, n196, n289, n290, n291, n749, n751, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788;
  wire   [287:0] STATE;

  OAI212 U3 ( .A(n289), .B(n1), .C(n293), .Q(n463) );
  OAI212 U5 ( .A(n289), .B(n2), .C(n295), .Q(n464) );
  OAI212 U7 ( .A(n289), .B(n3), .C(n296), .Q(n465) );
  OAI222 U9 ( .A(n196), .B(n3), .C(n773), .D(n4), .Q(n466) );
  OAI222 U10 ( .A(n757), .B(n4), .C(n771), .D(n5), .Q(n467) );
  OAI222 U11 ( .A(n760), .B(n5), .C(n772), .D(n6), .Q(n468) );
  OAI222 U12 ( .A(n764), .B(n6), .C(n774), .D(n7), .Q(n469) );
  OAI222 U13 ( .A(n763), .B(n7), .C(n772), .D(n8), .Q(n470) );
  OAI222 U14 ( .A(n760), .B(n8), .C(n771), .D(n9), .Q(n471) );
  OAI222 U15 ( .A(n758), .B(n9), .C(n771), .D(n10), .Q(n472) );
  OAI222 U16 ( .A(n760), .B(n10), .C(n769), .D(n11), .Q(n473) );
  OAI222 U17 ( .A(n749), .B(n11), .C(n774), .D(n12), .Q(n474) );
  OAI222 U18 ( .A(n758), .B(n12), .C(n770), .D(n13), .Q(n475) );
  OAI222 U19 ( .A(n196), .B(n13), .C(n775), .D(n14), .Q(n476) );
  OAI222 U20 ( .A(n758), .B(n14), .C(n775), .D(n15), .Q(n477) );
  OAI222 U21 ( .A(n757), .B(n15), .C(n775), .D(n16), .Q(n478) );
  OAI222 U22 ( .A(n757), .B(n16), .C(n775), .D(n17), .Q(n479) );
  OAI222 U23 ( .A(n757), .B(n17), .C(n775), .D(n18), .Q(n480) );
  OAI222 U24 ( .A(n757), .B(n18), .C(n775), .D(n19), .Q(n481) );
  OAI222 U25 ( .A(n757), .B(n19), .C(n775), .D(n20), .Q(n482) );
  OAI222 U26 ( .A(n757), .B(n20), .C(n774), .D(n21), .Q(n483) );
  OAI222 U27 ( .A(n757), .B(n21), .C(n774), .D(n22), .Q(n484) );
  OAI222 U28 ( .A(n757), .B(n22), .C(n774), .D(n23), .Q(n485) );
  OAI222 U29 ( .A(n757), .B(n23), .C(n774), .D(n24), .Q(n486) );
  OAI222 U30 ( .A(n757), .B(n24), .C(n774), .D(n26), .Q(n487) );
  OAI222 U31 ( .A(n757), .B(n26), .C(n774), .D(n27), .Q(n488) );
  OAI222 U32 ( .A(n757), .B(n27), .C(n774), .D(n28), .Q(n489) );
  OAI222 U33 ( .A(n757), .B(n28), .C(n775), .D(n29), .Q(n490) );
  OAI222 U34 ( .A(n749), .B(n29), .C(n770), .D(n30), .Q(n491) );
  OAI222 U35 ( .A(n757), .B(n30), .C(n770), .D(n31), .Q(n492) );
  OAI222 U36 ( .A(n196), .B(n31), .C(n775), .D(n32), .Q(n493) );
  OAI222 U37 ( .A(n758), .B(n32), .C(n773), .D(n33), .Q(n494) );
  OAI222 U38 ( .A(n196), .B(n33), .C(n772), .D(n34), .Q(n495) );
  OAI222 U39 ( .A(n196), .B(n34), .C(n769), .D(n35), .Q(n496) );
  OAI222 U40 ( .A(n749), .B(n35), .C(n772), .D(n36), .Q(n497) );
  OAI222 U41 ( .A(n756), .B(n36), .C(n771), .D(n37), .Q(n498) );
  OAI222 U42 ( .A(n763), .B(n37), .C(n770), .D(n38), .Q(n499) );
  OAI222 U43 ( .A(n756), .B(n38), .C(n775), .D(n39), .Q(n500) );
  OAI222 U44 ( .A(n764), .B(n39), .C(n770), .D(n40), .Q(n501) );
  OAI222 U45 ( .A(n749), .B(n40), .C(n773), .D(n41), .Q(n502) );
  OAI222 U46 ( .A(n762), .B(n41), .C(n775), .D(n42), .Q(n503) );
  OAI222 U47 ( .A(n757), .B(n42), .C(n773), .D(n43), .Q(n504) );
  OAI222 U48 ( .A(n196), .B(n43), .C(n773), .D(n44), .Q(n505) );
  OAI222 U49 ( .A(n758), .B(n44), .C(n773), .D(n45), .Q(n506) );
  OAI222 U50 ( .A(n751), .B(n45), .C(n773), .D(n46), .Q(n507) );
  OAI222 U51 ( .A(n757), .B(n46), .C(n773), .D(n47), .Q(n508) );
  OAI222 U52 ( .A(n751), .B(n47), .C(n773), .D(n48), .Q(n509) );
  OAI222 U53 ( .A(n749), .B(n48), .C(n773), .D(n49), .Q(n510) );
  OAI222 U54 ( .A(n756), .B(n49), .C(n771), .D(n50), .Q(n511) );
  OAI222 U55 ( .A(n762), .B(n50), .C(n769), .D(n51), .Q(n512) );
  OAI222 U56 ( .A(n761), .B(n51), .C(n774), .D(n52), .Q(n513) );
  OAI222 U57 ( .A(n760), .B(n52), .C(n776), .D(n53), .Q(n514) );
  OAI222 U58 ( .A(n749), .B(n53), .C(n772), .D(n54), .Q(n515) );
  OAI222 U59 ( .A(n749), .B(n54), .C(n771), .D(n55), .Q(n516) );
  OAI222 U60 ( .A(n751), .B(n55), .C(n769), .D(n56), .Q(n517) );
  OAI222 U61 ( .A(n759), .B(n56), .C(n769), .D(n57), .Q(n518) );
  OAI222 U62 ( .A(n757), .B(n57), .C(n771), .D(n58), .Q(n519) );
  OAI222 U63 ( .A(n757), .B(n58), .C(n773), .D(n59), .Q(n520) );
  OAI222 U64 ( .A(n196), .B(n59), .C(n770), .D(n60), .Q(n521) );
  OAI222 U65 ( .A(n196), .B(n60), .C(n774), .D(n61), .Q(n522) );
  OAI222 U66 ( .A(n196), .B(n61), .C(n769), .D(n62), .Q(n523) );
  OAI222 U67 ( .A(n196), .B(n62), .C(n774), .D(n63), .Q(n524) );
  OAI222 U68 ( .A(n196), .B(n63), .C(n771), .D(n64), .Q(n525) );
  OAI222 U69 ( .A(n749), .B(n64), .C(n771), .D(n65), .Q(n526) );
  OAI222 U70 ( .A(n751), .B(n65), .C(n769), .D(n66), .Q(n527) );
  OAI222 U71 ( .A(n756), .B(n66), .C(n774), .D(n67), .Q(n528) );
  OAI222 U72 ( .A(n759), .B(n67), .C(n772), .D(n68), .Q(n529) );
  OAI222 U73 ( .A(n196), .B(n68), .C(n770), .D(n69), .Q(n530) );
  OAI222 U74 ( .A(n758), .B(n69), .C(n775), .D(n70), .Q(n531) );
  OAI222 U75 ( .A(n764), .B(n70), .C(n772), .D(n71), .Q(n532) );
  OAI222 U76 ( .A(n749), .B(n71), .C(n772), .D(n72), .Q(n533) );
  OAI222 U77 ( .A(n751), .B(n72), .C(n772), .D(n73), .Q(n534) );
  OAI222 U78 ( .A(n756), .B(n73), .C(n772), .D(n74), .Q(n535) );
  OAI222 U79 ( .A(n751), .B(n74), .C(n772), .D(n75), .Q(n536) );
  OAI222 U80 ( .A(n196), .B(n75), .C(n772), .D(n76), .Q(n537) );
  OAI222 U81 ( .A(n196), .B(n76), .C(n772), .D(n77), .Q(n538) );
  OAI222 U82 ( .A(n758), .B(n77), .C(n771), .D(n78), .Q(n539) );
  OAI222 U83 ( .A(n749), .B(n78), .C(n771), .D(n79), .Q(n540) );
  OAI222 U84 ( .A(n756), .B(n79), .C(n771), .D(n80), .Q(n541) );
  OAI222 U85 ( .A(n751), .B(n80), .C(n771), .D(n81), .Q(n542) );
  OAI222 U86 ( .A(n196), .B(n81), .C(n771), .D(n82), .Q(n543) );
  OAI222 U87 ( .A(n196), .B(n82), .C(n771), .D(n83), .Q(n544) );
  OAI222 U88 ( .A(n758), .B(n83), .C(n771), .D(n84), .Q(n545) );
  OAI222 U89 ( .A(n749), .B(n84), .C(n775), .D(n85), .Q(n546) );
  OAI222 U90 ( .A(n756), .B(n85), .C(n773), .D(n86), .Q(n547) );
  OAI222 U91 ( .A(n751), .B(n86), .C(n776), .D(n87), .Q(n548) );
  OAI222 U92 ( .A(n196), .B(n87), .C(n769), .D(n88), .Q(n549) );
  OAI222 U93 ( .A(n763), .B(n88), .C(n774), .D(n89), .Q(n550) );
  OAI222 U94 ( .A(n763), .B(n89), .C(n772), .D(n90), .Q(n551) );
  OAI222 U95 ( .A(n763), .B(n90), .C(n771), .D(n91), .Q(n552) );
  OAI222 U96 ( .A(n763), .B(n91), .C(n772), .D(n92), .Q(n553) );
  OAI222 U97 ( .A(n763), .B(n92), .C(n776), .D(n93), .Q(n554) );
  OAI222 U98 ( .A(n763), .B(n93), .C(n769), .D(n94), .Q(n555) );
  OAI222 U99 ( .A(n763), .B(n94), .C(n774), .D(n95), .Q(n556) );
  OAI222 U100 ( .A(n763), .B(n95), .C(n772), .D(n96), .Q(n557) );
  OAI222 U101 ( .A(n763), .B(n96), .C(n771), .D(n97), .Q(n558) );
  OAI222 U102 ( .A(n763), .B(n97), .C(n776), .D(n98), .Q(n559) );
  OAI222 U103 ( .A(n763), .B(n98), .C(n770), .D(n99), .Q(n560) );
  OAI222 U104 ( .A(n763), .B(n99), .C(n770), .D(n100), .Q(n561) );
  OAI222 U105 ( .A(n763), .B(n100), .C(n770), .D(n101), .Q(n562) );
  OAI222 U106 ( .A(n763), .B(n101), .C(n770), .D(n102), .Q(n563) );
  OAI222 U107 ( .A(n763), .B(n102), .C(n770), .D(n103), .Q(n564) );
  OAI222 U108 ( .A(n764), .B(n103), .C(n770), .D(n104), .Q(n565) );
  OAI222 U109 ( .A(n764), .B(n104), .C(n770), .D(n105), .Q(n566) );
  OAI222 U110 ( .A(n764), .B(n105), .C(n769), .D(n106), .Q(n567) );
  OAI222 U111 ( .A(n764), .B(n106), .C(n769), .D(n107), .Q(n568) );
  OAI222 U112 ( .A(n764), .B(n107), .C(n769), .D(n108), .Q(n569) );
  OAI222 U113 ( .A(n764), .B(n108), .C(n769), .D(n109), .Q(n570) );
  OAI222 U118 ( .A(n764), .B(n113), .C(n769), .D(n114), .Q(n571) );
  OAI222 U119 ( .A(n764), .B(n114), .C(n769), .D(n115), .Q(n572) );
  OAI222 U120 ( .A(n764), .B(n115), .C(n769), .D(n116), .Q(n573) );
  OAI212 U121 ( .A(n751), .B(n116), .C(n302), .Q(n574) );
  OAI212 U123 ( .A(n758), .B(n117), .C(n303), .Q(n575) );
  OAI212 U125 ( .A(n758), .B(n118), .C(n304), .Q(n576) );
  OAI212 U127 ( .A(n763), .B(n119), .C(n305), .Q(n577) );
  OAI212 U129 ( .A(n760), .B(n120), .C(n306), .Q(n578) );
  OAI212 U131 ( .A(n763), .B(n121), .C(n307), .Q(n579) );
  OAI212 U133 ( .A(n759), .B(n122), .C(n308), .Q(n580) );
  OAI212 U135 ( .A(n757), .B(n123), .C(n309), .Q(n581) );
  OAI212 U137 ( .A(n758), .B(n124), .C(n310), .Q(n582) );
  OAI212 U139 ( .A(n764), .B(n125), .C(n311), .Q(n583) );
  OAI212 U141 ( .A(n764), .B(n126), .C(n312), .Q(n584) );
  OAI212 U143 ( .A(n764), .B(n127), .C(n313), .Q(n585) );
  OAI212 U145 ( .A(n759), .B(n128), .C(n314), .Q(n586) );
  OAI212 U147 ( .A(n751), .B(n129), .C(n315), .Q(n587) );
  OAI212 U149 ( .A(n749), .B(n130), .C(n316), .Q(n588) );
  OAI212 U151 ( .A(n756), .B(n131), .C(n317), .Q(n589) );
  OAI212 U153 ( .A(n196), .B(n132), .C(n318), .Q(n590) );
  OAI212 U155 ( .A(n756), .B(n133), .C(n319), .Q(n591) );
  OAI212 U157 ( .A(n760), .B(n134), .C(n320), .Q(n592) );
  OAI212 U159 ( .A(n749), .B(n135), .C(n321), .Q(n593) );
  OAI212 U161 ( .A(n758), .B(n136), .C(n322), .Q(n594) );
  OAI212 U163 ( .A(n764), .B(n137), .C(n323), .Q(n595) );
  OAI212 U165 ( .A(n757), .B(n138), .C(n324), .Q(n596) );
  OAI212 U167 ( .A(n751), .B(n139), .C(n325), .Q(n597) );
  OAI212 U169 ( .A(n762), .B(n140), .C(n326), .Q(n598) );
  OAI212 U171 ( .A(n761), .B(n141), .C(n327), .Q(n599) );
  OAI212 U173 ( .A(n196), .B(n142), .C(n328), .Q(n600) );
  OAI212 U175 ( .A(n751), .B(n143), .C(n329), .Q(n601) );
  OAI212 U177 ( .A(n196), .B(n144), .C(n330), .Q(n602) );
  OAI212 U179 ( .A(n749), .B(n145), .C(n331), .Q(n603) );
  OAI212 U181 ( .A(n758), .B(n146), .C(n332), .Q(n604) );
  OAI212 U183 ( .A(n763), .B(n147), .C(n333), .Q(n605) );
  OAI212 U185 ( .A(n756), .B(n148), .C(n334), .Q(n606) );
  OAI212 U187 ( .A(n757), .B(n149), .C(n335), .Q(n607) );
  OAI212 U189 ( .A(n756), .B(n150), .C(n336), .Q(n608) );
  OAI212 U191 ( .A(n196), .B(n151), .C(n337), .Q(n609) );
  OAI212 U193 ( .A(n759), .B(n152), .C(n338), .Q(n610) );
  OAI212 U195 ( .A(n196), .B(n153), .C(n339), .Q(n611) );
  OAI212 U197 ( .A(n751), .B(n154), .C(n340), .Q(n612) );
  OAI212 U199 ( .A(n759), .B(n155), .C(n341), .Q(n613) );
  OAI212 U201 ( .A(n751), .B(n156), .C(n342), .Q(n614) );
  OAI212 U203 ( .A(n749), .B(n157), .C(n343), .Q(n615) );
  OAI212 U205 ( .A(n760), .B(n158), .C(n344), .Q(n616) );
  OAI212 U207 ( .A(n762), .B(n159), .C(n345), .Q(n617) );
  OAI212 U209 ( .A(n751), .B(n160), .C(n346), .Q(n618) );
  OAI212 U211 ( .A(n758), .B(n161), .C(n347), .Q(n619) );
  OAI212 U213 ( .A(n763), .B(n162), .C(n348), .Q(n620) );
  OAI212 U215 ( .A(n756), .B(n163), .C(n349), .Q(n621) );
  OAI212 U217 ( .A(n763), .B(n164), .C(n350), .Q(n622) );
  OAI212 U219 ( .A(n751), .B(n165), .C(n351), .Q(n623) );
  OAI212 U221 ( .A(n196), .B(n166), .C(n352), .Q(n624) );
  OAI212 U223 ( .A(n759), .B(n167), .C(n353), .Q(n625) );
  OAI212 U225 ( .A(n764), .B(n168), .C(n354), .Q(n626) );
  OAI212 U227 ( .A(n196), .B(n169), .C(n355), .Q(n627) );
  OAI212 U229 ( .A(n751), .B(n170), .C(n356), .Q(n628) );
  OAI212 U231 ( .A(n763), .B(n171), .C(n357), .Q(n629) );
  OAI212 U233 ( .A(n749), .B(n172), .C(n358), .Q(n630) );
  OAI212 U235 ( .A(n756), .B(n173), .C(n359), .Q(n631) );
  OAI212 U237 ( .A(n764), .B(n174), .C(n360), .Q(n632) );
  OAI212 U239 ( .A(n763), .B(n175), .C(n361), .Q(n633) );
  OAI212 U241 ( .A(n196), .B(n176), .C(n362), .Q(n634) );
  OAI212 U243 ( .A(n751), .B(n177), .C(n363), .Q(n635) );
  OAI212 U245 ( .A(n762), .B(n178), .C(n364), .Q(n636) );
  OAI212 U247 ( .A(n761), .B(n179), .C(n365), .Q(n637) );
  OAI212 U249 ( .A(n749), .B(n180), .C(n366), .Q(n638) );
  OAI212 U251 ( .A(n759), .B(n181), .C(n367), .Q(n639) );
  OAI212 U253 ( .A(n759), .B(n182), .C(n368), .Q(n640) );
  OAI212 U255 ( .A(n759), .B(n183), .C(n369), .Q(n641) );
  OAI212 U257 ( .A(n759), .B(n184), .C(n370), .Q(n642) );
  OAI212 U259 ( .A(n759), .B(n185), .C(n371), .Q(n643) );
  OAI212 U261 ( .A(n759), .B(n186), .C(n372), .Q(n644) );
  OAI212 U263 ( .A(n759), .B(n187), .C(n373), .Q(n645) );
  OAI212 U265 ( .A(n759), .B(n188), .C(n374), .Q(n646) );
  OAI212 U267 ( .A(n759), .B(n189), .C(n375), .Q(n647) );
  OAI212 U269 ( .A(n759), .B(n190), .C(n376), .Q(n648) );
  OAI212 U271 ( .A(n759), .B(n191), .C(n377), .Q(n649) );
  OAI212 U273 ( .A(n759), .B(n192), .C(n378), .Q(n650) );
  OAI212 U275 ( .A(n759), .B(n193), .C(n379), .Q(n651) );
  OAI212 U277 ( .A(n760), .B(n194), .C(n380), .Q(n652) );
  OAI212 U279 ( .A(n760), .B(n195), .C(n381), .Q(n653) );
  OAI222 U282 ( .A(n764), .B(n197), .C(n770), .D(n198), .Q(n654) );
  OAI222 U283 ( .A(n764), .B(n198), .C(n775), .D(n199), .Q(n655) );
  OAI222 U284 ( .A(n764), .B(n199), .C(n773), .D(n200), .Q(n656) );
  OAI222 U285 ( .A(n764), .B(n200), .C(n773), .D(n201), .Q(n657) );
  OAI222 U286 ( .A(n764), .B(n201), .C(n769), .D(n202), .Q(n658) );
  OAI222 U287 ( .A(n763), .B(n202), .C(n774), .D(n203), .Q(n659) );
  OAI222 U288 ( .A(n196), .B(n203), .C(n772), .D(n204), .Q(n660) );
  OAI222 U289 ( .A(n749), .B(n204), .C(n773), .D(n205), .Q(n661) );
  OAI222 U290 ( .A(n757), .B(n205), .C(n775), .D(n206), .Q(n662) );
  OAI222 U291 ( .A(n759), .B(n206), .C(n769), .D(n207), .Q(n663) );
  OAI222 U292 ( .A(n757), .B(n207), .C(n774), .D(n208), .Q(n664) );
  OAI222 U293 ( .A(n764), .B(n208), .C(n772), .D(n209), .Q(n665) );
  OAI212 U294 ( .A(n757), .B(n209), .C(n383), .Q(n666) );
  OAI212 U296 ( .A(n764), .B(n210), .C(n384), .Q(n667) );
  OAI212 U298 ( .A(n757), .B(n211), .C(n385), .Q(n668) );
  OAI212 U300 ( .A(n760), .B(n212), .C(n386), .Q(n669) );
  OAI212 U302 ( .A(n760), .B(n213), .C(n387), .Q(n670) );
  OAI212 U304 ( .A(n758), .B(n214), .C(n388), .Q(n671) );
  OAI212 U306 ( .A(n756), .B(n215), .C(n389), .Q(n672) );
  OAI212 U308 ( .A(n756), .B(n216), .C(n390), .Q(n673) );
  OAI212 U310 ( .A(n749), .B(n217), .C(n391), .Q(n674) );
  OAI212 U312 ( .A(n751), .B(n218), .C(n392), .Q(n675) );
  OAI212 U314 ( .A(n758), .B(n219), .C(n393), .Q(n676) );
  OAI212 U316 ( .A(n756), .B(n220), .C(n394), .Q(n677) );
  OAI212 U318 ( .A(n749), .B(n221), .C(n395), .Q(n678) );
  OAI212 U320 ( .A(n751), .B(n222), .C(n396), .Q(n679) );
  OAI212 U322 ( .A(n758), .B(n223), .C(n397), .Q(n680) );
  OAI212 U324 ( .A(n756), .B(n224), .C(n398), .Q(n681) );
  OAI212 U326 ( .A(n749), .B(n225), .C(n399), .Q(n682) );
  OAI212 U328 ( .A(n751), .B(n226), .C(n400), .Q(n683) );
  OAI212 U330 ( .A(n751), .B(n227), .C(n401), .Q(n684) );
  OAI212 U332 ( .A(n759), .B(n228), .C(n402), .Q(n685) );
  OAI212 U334 ( .A(n756), .B(n229), .C(n403), .Q(n686) );
  OAI212 U336 ( .A(n758), .B(n230), .C(n404), .Q(n687) );
  OAI212 U338 ( .A(n196), .B(n231), .C(n405), .Q(n688) );
  OAI212 U340 ( .A(n196), .B(n232), .C(n406), .Q(n689) );
  OAI212 U342 ( .A(n196), .B(n233), .C(n407), .Q(n690) );
  OAI212 U344 ( .A(n196), .B(n234), .C(n408), .Q(n691) );
  OAI212 U346 ( .A(n196), .B(n235), .C(n409), .Q(n692) );
  OAI212 U348 ( .A(n196), .B(n236), .C(n410), .Q(n693) );
  OAI212 U350 ( .A(n196), .B(n237), .C(n411), .Q(n694) );
  OAI212 U352 ( .A(n761), .B(n238), .C(n412), .Q(n695) );
  OAI212 U354 ( .A(n762), .B(n239), .C(n413), .Q(n696) );
  OAI212 U356 ( .A(n762), .B(n240), .C(n414), .Q(n697) );
  OAI212 U358 ( .A(n762), .B(n241), .C(n415), .Q(n698) );
  OAI212 U360 ( .A(n762), .B(n242), .C(n416), .Q(n699) );
  OAI212 U362 ( .A(n762), .B(n243), .C(n417), .Q(n700) );
  OAI212 U364 ( .A(n762), .B(n244), .C(n418), .Q(n701) );
  OAI212 U366 ( .A(n762), .B(n245), .C(n419), .Q(n702) );
  OAI212 U368 ( .A(n762), .B(n246), .C(n420), .Q(n703) );
  OAI212 U370 ( .A(n762), .B(n247), .C(n421), .Q(n704) );
  OAI212 U372 ( .A(n762), .B(n248), .C(n422), .Q(n705) );
  OAI212 U374 ( .A(n762), .B(n249), .C(n423), .Q(n706) );
  OAI212 U376 ( .A(n762), .B(n250), .C(n424), .Q(n707) );
  OAI212 U378 ( .A(n761), .B(n251), .C(n425), .Q(n708) );
  OAI212 U380 ( .A(n761), .B(n252), .C(n426), .Q(n709) );
  OAI212 U382 ( .A(n761), .B(n253), .C(n427), .Q(n710) );
  OAI212 U384 ( .A(n761), .B(n254), .C(n428), .Q(n711) );
  OAI212 U386 ( .A(n761), .B(n255), .C(n429), .Q(n712) );
  OAI212 U388 ( .A(n761), .B(n256), .C(n430), .Q(n713) );
  OAI212 U390 ( .A(n761), .B(n257), .C(n431), .Q(n714) );
  OAI212 U392 ( .A(n761), .B(n258), .C(n432), .Q(n715) );
  OAI212 U394 ( .A(n761), .B(n259), .C(n433), .Q(n716) );
  OAI212 U396 ( .A(n761), .B(n260), .C(n434), .Q(n717) );
  OAI212 U398 ( .A(n761), .B(n261), .C(n435), .Q(n718) );
  OAI212 U400 ( .A(n761), .B(n262), .C(n436), .Q(n719) );
  OAI212 U402 ( .A(n761), .B(n263), .C(n437), .Q(n720) );
  OAI212 U404 ( .A(n758), .B(n264), .C(n438), .Q(n721) );
  OAI212 U406 ( .A(n756), .B(n265), .C(n439), .Q(n722) );
  OAI212 U408 ( .A(n761), .B(n266), .C(n440), .Q(n723) );
  OAI212 U410 ( .A(n762), .B(n267), .C(n441), .Q(n724) );
  OAI212 U412 ( .A(n749), .B(n268), .C(n442), .Q(n725) );
  OAI212 U414 ( .A(n758), .B(n269), .C(n443), .Q(n726) );
  OAI212 U416 ( .A(n756), .B(n270), .C(n444), .Q(n727) );
  OAI212 U418 ( .A(n761), .B(n271), .C(n445), .Q(n728) );
  OAI212 U420 ( .A(n762), .B(n272), .C(n446), .Q(n729) );
  OAI212 U422 ( .A(n749), .B(n273), .C(n447), .Q(n730) );
  OAI212 U424 ( .A(n758), .B(n274), .C(n448), .Q(n731) );
  OAI212 U426 ( .A(n756), .B(n275), .C(n449), .Q(n732) );
  OAI212 U428 ( .A(n761), .B(n276), .C(n450), .Q(n733) );
  OAI212 U430 ( .A(n760), .B(n277), .C(n451), .Q(n734) );
  OAI212 U432 ( .A(n760), .B(n278), .C(n452), .Q(n735) );
  OAI212 U434 ( .A(n760), .B(n279), .C(n453), .Q(n736) );
  OAI212 U436 ( .A(n760), .B(n280), .C(n454), .Q(n737) );
  OAI212 U438 ( .A(n760), .B(n281), .C(n455), .Q(n738) );
  OAI212 U440 ( .A(n760), .B(n282), .C(n456), .Q(n739) );
  OAI212 U442 ( .A(n760), .B(n283), .C(n457), .Q(n740) );
  OAI212 U444 ( .A(n760), .B(n284), .C(n458), .Q(n741) );
  OAI212 U446 ( .A(n760), .B(n285), .C(n459), .Q(n742) );
  OAI212 U448 ( .A(n760), .B(n286), .C(n460), .Q(n743) );
  OAI212 U450 ( .A(n760), .B(n287), .C(n461), .Q(n744) );
  OAI212 U452 ( .A(n762), .B(n288), .C(n462), .Q(n745) );
  DF3 STATE_reg_0_ ( .D(n745), .C(SYS_CLK), .Q(STATE[0]), .QN(n288) );
  DF3 STATE_reg_1_ ( .D(n744), .C(SYS_CLK), .Q(STATE[1]), .QN(n287) );
  DF3 STATE_reg_2_ ( .D(n743), .C(SYS_CLK), .Q(STATE[2]), .QN(n286) );
  DF3 STATE_reg_3_ ( .D(n742), .C(SYS_CLK), .Q(STATE[3]), .QN(n285) );
  DF3 STATE_reg_4_ ( .D(n741), .C(SYS_CLK), .Q(STATE[4]), .QN(n284) );
  DF3 STATE_reg_5_ ( .D(n740), .C(SYS_CLK), .Q(STATE[5]), .QN(n283) );
  DF3 STATE_reg_6_ ( .D(n739), .C(SYS_CLK), .Q(STATE[6]), .QN(n282) );
  DF3 STATE_reg_7_ ( .D(n738), .C(SYS_CLK), .Q(STATE[7]), .QN(n281) );
  DF3 STATE_reg_8_ ( .D(n737), .C(SYS_CLK), .Q(STATE[8]), .QN(n280) );
  DF3 STATE_reg_9_ ( .D(n736), .C(SYS_CLK), .Q(STATE[9]), .QN(n279) );
  DF3 STATE_reg_10_ ( .D(n735), .C(SYS_CLK), .Q(STATE[10]), .QN(n278) );
  DF3 STATE_reg_11_ ( .D(n734), .C(SYS_CLK), .Q(STATE[11]), .QN(n277) );
  DF3 STATE_reg_12_ ( .D(n733), .C(SYS_CLK), .Q(STATE[12]), .QN(n276) );
  DF3 STATE_reg_13_ ( .D(n732), .C(SYS_CLK), .Q(STATE[13]), .QN(n275) );
  DF3 STATE_reg_14_ ( .D(n731), .C(SYS_CLK), .Q(STATE[14]), .QN(n274) );
  DF3 STATE_reg_15_ ( .D(n730), .C(SYS_CLK), .Q(STATE[15]), .QN(n273) );
  DF3 STATE_reg_16_ ( .D(n729), .C(SYS_CLK), .Q(STATE[16]), .QN(n272) );
  DF3 STATE_reg_17_ ( .D(n728), .C(SYS_CLK), .Q(STATE[17]), .QN(n271) );
  DF3 STATE_reg_18_ ( .D(n727), .C(SYS_CLK), .Q(STATE[18]), .QN(n270) );
  DF3 STATE_reg_19_ ( .D(n726), .C(SYS_CLK), .Q(STATE[19]), .QN(n269) );
  DF3 STATE_reg_20_ ( .D(n725), .C(SYS_CLK), .Q(STATE[20]), .QN(n268) );
  DF3 STATE_reg_21_ ( .D(n724), .C(SYS_CLK), .Q(STATE[21]), .QN(n267) );
  DF3 STATE_reg_22_ ( .D(n723), .C(SYS_CLK), .Q(STATE[22]), .QN(n266) );
  DF3 STATE_reg_23_ ( .D(n722), .C(SYS_CLK), .Q(STATE[23]), .QN(n265) );
  DF3 STATE_reg_24_ ( .D(n721), .C(SYS_CLK), .Q(STATE[24]), .QN(n264) );
  DF3 STATE_reg_25_ ( .D(n720), .C(SYS_CLK), .Q(STATE[25]), .QN(n263) );
  DF3 STATE_reg_26_ ( .D(n719), .C(SYS_CLK), .Q(STATE[26]), .QN(n262) );
  DF3 STATE_reg_27_ ( .D(n718), .C(SYS_CLK), .Q(STATE[27]), .QN(n261) );
  DF3 STATE_reg_28_ ( .D(n717), .C(SYS_CLK), .Q(STATE[28]), .QN(n260) );
  DF3 STATE_reg_29_ ( .D(n716), .C(SYS_CLK), .Q(STATE[29]), .QN(n259) );
  DF3 STATE_reg_30_ ( .D(n715), .C(SYS_CLK), .Q(STATE[30]), .QN(n258) );
  DF3 STATE_reg_31_ ( .D(n714), .C(SYS_CLK), .Q(STATE[31]), .QN(n257) );
  DF3 STATE_reg_32_ ( .D(n713), .C(SYS_CLK), .Q(STATE[32]), .QN(n256) );
  DF3 STATE_reg_33_ ( .D(n712), .C(SYS_CLK), .Q(STATE[33]), .QN(n255) );
  DF3 STATE_reg_34_ ( .D(n711), .C(SYS_CLK), .Q(STATE[34]), .QN(n254) );
  DF3 STATE_reg_35_ ( .D(n710), .C(SYS_CLK), .Q(STATE[35]), .QN(n253) );
  DF3 STATE_reg_36_ ( .D(n709), .C(SYS_CLK), .Q(STATE[36]), .QN(n252) );
  DF3 STATE_reg_37_ ( .D(n708), .C(SYS_CLK), .Q(STATE[37]), .QN(n251) );
  DF3 STATE_reg_38_ ( .D(n707), .C(SYS_CLK), .Q(STATE[38]), .QN(n250) );
  DF3 STATE_reg_39_ ( .D(n706), .C(SYS_CLK), .Q(STATE[39]), .QN(n249) );
  DF3 STATE_reg_40_ ( .D(n705), .C(SYS_CLK), .Q(STATE[40]), .QN(n248) );
  DF3 STATE_reg_41_ ( .D(n704), .C(SYS_CLK), .Q(STATE[41]), .QN(n247) );
  DF3 STATE_reg_42_ ( .D(n703), .C(SYS_CLK), .Q(STATE[42]), .QN(n246) );
  DF3 STATE_reg_43_ ( .D(n702), .C(SYS_CLK), .Q(STATE[43]), .QN(n245) );
  DF3 STATE_reg_44_ ( .D(n701), .C(SYS_CLK), .Q(STATE[44]), .QN(n244) );
  DF3 STATE_reg_45_ ( .D(n700), .C(SYS_CLK), .Q(STATE[45]), .QN(n243) );
  DF3 STATE_reg_46_ ( .D(n699), .C(SYS_CLK), .Q(STATE[46]), .QN(n242) );
  DF3 STATE_reg_47_ ( .D(n698), .C(SYS_CLK), .Q(STATE[47]), .QN(n241) );
  DF3 STATE_reg_48_ ( .D(n697), .C(SYS_CLK), .Q(STATE[48]), .QN(n240) );
  DF3 STATE_reg_49_ ( .D(n696), .C(SYS_CLK), .Q(STATE[49]), .QN(n239) );
  DF3 STATE_reg_50_ ( .D(n695), .C(SYS_CLK), .Q(STATE[50]), .QN(n238) );
  DF3 STATE_reg_51_ ( .D(n694), .C(SYS_CLK), .Q(STATE[51]), .QN(n237) );
  DF3 STATE_reg_52_ ( .D(n693), .C(SYS_CLK), .Q(STATE[52]), .QN(n236) );
  DF3 STATE_reg_53_ ( .D(n692), .C(SYS_CLK), .Q(STATE[53]), .QN(n235) );
  DF3 STATE_reg_54_ ( .D(n691), .C(SYS_CLK), .Q(STATE[54]), .QN(n234) );
  DF3 STATE_reg_55_ ( .D(n690), .C(SYS_CLK), .Q(STATE[55]), .QN(n233) );
  DF3 STATE_reg_56_ ( .D(n689), .C(SYS_CLK), .Q(STATE[56]), .QN(n232) );
  DF3 STATE_reg_57_ ( .D(n688), .C(SYS_CLK), .Q(STATE[57]), .QN(n231) );
  DF3 STATE_reg_58_ ( .D(n687), .C(SYS_CLK), .Q(STATE[58]), .QN(n230) );
  DF3 STATE_reg_59_ ( .D(n686), .C(SYS_CLK), .Q(STATE[59]), .QN(n229) );
  DF3 STATE_reg_60_ ( .D(n685), .C(SYS_CLK), .Q(STATE[60]), .QN(n228) );
  DF3 STATE_reg_61_ ( .D(n684), .C(SYS_CLK), .Q(STATE[61]), .QN(n227) );
  DF3 STATE_reg_62_ ( .D(n683), .C(SYS_CLK), .Q(STATE[62]), .QN(n226) );
  DF3 STATE_reg_63_ ( .D(n682), .C(SYS_CLK), .Q(STATE[63]), .QN(n225) );
  DF3 STATE_reg_64_ ( .D(n681), .C(SYS_CLK), .Q(STATE[64]), .QN(n224) );
  DF3 STATE_reg_65_ ( .D(n680), .C(SYS_CLK), .Q(STATE[65]), .QN(n223) );
  DF3 STATE_reg_66_ ( .D(n679), .C(SYS_CLK), .Q(STATE[66]), .QN(n222) );
  DF3 STATE_reg_67_ ( .D(n678), .C(SYS_CLK), .Q(STATE[67]), .QN(n221) );
  DF3 STATE_reg_68_ ( .D(n677), .C(SYS_CLK), .Q(STATE[68]), .QN(n220) );
  DF3 STATE_reg_69_ ( .D(n676), .C(SYS_CLK), .Q(STATE[69]), .QN(n219) );
  DF3 STATE_reg_70_ ( .D(n675), .C(SYS_CLK), .Q(STATE[70]), .QN(n218) );
  DF3 STATE_reg_71_ ( .D(n674), .C(SYS_CLK), .Q(STATE[71]), .QN(n217) );
  DF3 STATE_reg_72_ ( .D(n673), .C(SYS_CLK), .Q(STATE[72]), .QN(n216) );
  DF3 STATE_reg_73_ ( .D(n672), .C(SYS_CLK), .Q(STATE[73]), .QN(n215) );
  DF3 STATE_reg_74_ ( .D(n671), .C(SYS_CLK), .Q(STATE[74]), .QN(n214) );
  DF3 STATE_reg_75_ ( .D(n670), .C(SYS_CLK), .Q(STATE[75]), .QN(n213) );
  DF3 STATE_reg_76_ ( .D(n669), .C(SYS_CLK), .Q(STATE[76]), .QN(n212) );
  DF3 STATE_reg_77_ ( .D(n668), .C(SYS_CLK), .Q(STATE[77]), .QN(n211) );
  DF3 STATE_reg_78_ ( .D(n667), .C(SYS_CLK), .Q(STATE[78]), .QN(n210) );
  DF3 STATE_reg_79_ ( .D(n666), .C(SYS_CLK), .QN(n209) );
  DF3 STATE_reg_80_ ( .D(n665), .C(SYS_CLK), .QN(n208) );
  DF3 STATE_reg_81_ ( .D(n664), .C(SYS_CLK), .QN(n207) );
  DF3 STATE_reg_82_ ( .D(n663), .C(SYS_CLK), .QN(n206) );
  DF3 STATE_reg_83_ ( .D(n662), .C(SYS_CLK), .QN(n205) );
  DF3 STATE_reg_84_ ( .D(n661), .C(SYS_CLK), .QN(n204) );
  DF3 STATE_reg_85_ ( .D(n660), .C(SYS_CLK), .QN(n203) );
  DF3 STATE_reg_86_ ( .D(n659), .C(SYS_CLK), .QN(n202) );
  DF3 STATE_reg_87_ ( .D(n658), .C(SYS_CLK), .QN(n201) );
  DF3 STATE_reg_88_ ( .D(n657), .C(SYS_CLK), .QN(n200) );
  DF3 STATE_reg_89_ ( .D(n656), .C(SYS_CLK), .QN(n199) );
  DF3 STATE_reg_90_ ( .D(n655), .C(SYS_CLK), .QN(n198) );
  DF3 STATE_reg_91_ ( .D(n654), .C(SYS_CLK), .Q(STATE[91]), .QN(n197) );
  DF3 STATE_reg_92_ ( .D(n783), .C(SYS_CLK), .Q(STATE[92]) );
  DF3 STATE_reg_93_ ( .D(n653), .C(SYS_CLK), .Q(STATE[93]), .QN(n195) );
  DF3 STATE_reg_94_ ( .D(n652), .C(SYS_CLK), .Q(STATE[94]), .QN(n194) );
  DF3 STATE_reg_95_ ( .D(n651), .C(SYS_CLK), .Q(STATE[95]), .QN(n193) );
  DF3 STATE_reg_96_ ( .D(n650), .C(SYS_CLK), .Q(STATE[96]), .QN(n192) );
  DF3 STATE_reg_97_ ( .D(n649), .C(SYS_CLK), .Q(STATE[97]), .QN(n191) );
  DF3 STATE_reg_98_ ( .D(n648), .C(SYS_CLK), .Q(STATE[98]), .QN(n190) );
  DF3 STATE_reg_99_ ( .D(n647), .C(SYS_CLK), .Q(STATE[99]), .QN(n189) );
  DF3 STATE_reg_100_ ( .D(n646), .C(SYS_CLK), .Q(STATE[100]), .QN(n188) );
  DF3 STATE_reg_101_ ( .D(n645), .C(SYS_CLK), .Q(STATE[101]), .QN(n187) );
  DF3 STATE_reg_102_ ( .D(n644), .C(SYS_CLK), .Q(STATE[102]), .QN(n186) );
  DF3 STATE_reg_103_ ( .D(n643), .C(SYS_CLK), .Q(STATE[103]), .QN(n185) );
  DF3 STATE_reg_104_ ( .D(n642), .C(SYS_CLK), .Q(STATE[104]), .QN(n184) );
  DF3 STATE_reg_105_ ( .D(n641), .C(SYS_CLK), .Q(STATE[105]), .QN(n183) );
  DF3 STATE_reg_106_ ( .D(n640), .C(SYS_CLK), .Q(STATE[106]), .QN(n182) );
  DF3 STATE_reg_107_ ( .D(n639), .C(SYS_CLK), .Q(STATE[107]), .QN(n181) );
  DF3 STATE_reg_108_ ( .D(n638), .C(SYS_CLK), .Q(STATE[108]), .QN(n180) );
  DF3 STATE_reg_109_ ( .D(n637), .C(SYS_CLK), .Q(STATE[109]), .QN(n179) );
  DF3 STATE_reg_110_ ( .D(n636), .C(SYS_CLK), .Q(STATE[110]), .QN(n178) );
  DF3 STATE_reg_111_ ( .D(n635), .C(SYS_CLK), .Q(STATE[111]), .QN(n177) );
  DF3 STATE_reg_112_ ( .D(n634), .C(SYS_CLK), .Q(STATE[112]), .QN(n176) );
  DF3 STATE_reg_113_ ( .D(n633), .C(SYS_CLK), .Q(STATE[113]), .QN(n175) );
  DF3 STATE_reg_114_ ( .D(n632), .C(SYS_CLK), .Q(STATE[114]), .QN(n174) );
  DF3 STATE_reg_115_ ( .D(n631), .C(SYS_CLK), .Q(STATE[115]), .QN(n173) );
  DF3 STATE_reg_116_ ( .D(n630), .C(SYS_CLK), .Q(STATE[116]), .QN(n172) );
  DF3 STATE_reg_117_ ( .D(n629), .C(SYS_CLK), .Q(STATE[117]), .QN(n171) );
  DF3 STATE_reg_118_ ( .D(n628), .C(SYS_CLK), .Q(STATE[118]), .QN(n170) );
  DF3 STATE_reg_119_ ( .D(n627), .C(SYS_CLK), .Q(STATE[119]), .QN(n169) );
  DF3 STATE_reg_120_ ( .D(n626), .C(SYS_CLK), .Q(STATE[120]), .QN(n168) );
  DF3 STATE_reg_121_ ( .D(n625), .C(SYS_CLK), .Q(STATE[121]), .QN(n167) );
  DF3 STATE_reg_122_ ( .D(n624), .C(SYS_CLK), .Q(STATE[122]), .QN(n166) );
  DF3 STATE_reg_123_ ( .D(n623), .C(SYS_CLK), .Q(STATE[123]), .QN(n165) );
  DF3 STATE_reg_124_ ( .D(n622), .C(SYS_CLK), .Q(STATE[124]), .QN(n164) );
  DF3 STATE_reg_125_ ( .D(n621), .C(SYS_CLK), .Q(STATE[125]), .QN(n163) );
  DF3 STATE_reg_126_ ( .D(n620), .C(SYS_CLK), .Q(STATE[126]), .QN(n162) );
  DF3 STATE_reg_127_ ( .D(n619), .C(SYS_CLK), .Q(STATE[127]), .QN(n161) );
  DF3 STATE_reg_128_ ( .D(n618), .C(SYS_CLK), .Q(STATE[128]), .QN(n160) );
  DF3 STATE_reg_129_ ( .D(n617), .C(SYS_CLK), .Q(STATE[129]), .QN(n159) );
  DF3 STATE_reg_130_ ( .D(n616), .C(SYS_CLK), .Q(STATE[130]), .QN(n158) );
  DF3 STATE_reg_131_ ( .D(n615), .C(SYS_CLK), .Q(STATE[131]), .QN(n157) );
  DF3 STATE_reg_132_ ( .D(n614), .C(SYS_CLK), .Q(STATE[132]), .QN(n156) );
  DF3 STATE_reg_133_ ( .D(n613), .C(SYS_CLK), .Q(STATE[133]), .QN(n155) );
  DF3 STATE_reg_134_ ( .D(n612), .C(SYS_CLK), .Q(STATE[134]), .QN(n154) );
  DF3 STATE_reg_135_ ( .D(n611), .C(SYS_CLK), .Q(STATE[135]), .QN(n153) );
  DF3 STATE_reg_136_ ( .D(n610), .C(SYS_CLK), .Q(STATE[136]), .QN(n152) );
  DF3 STATE_reg_137_ ( .D(n609), .C(SYS_CLK), .Q(STATE[137]), .QN(n151) );
  DF3 STATE_reg_138_ ( .D(n608), .C(SYS_CLK), .Q(STATE[138]), .QN(n150) );
  DF3 STATE_reg_139_ ( .D(n607), .C(SYS_CLK), .Q(STATE[139]), .QN(n149) );
  DF3 STATE_reg_140_ ( .D(n606), .C(SYS_CLK), .Q(STATE[140]), .QN(n148) );
  DF3 STATE_reg_141_ ( .D(n605), .C(SYS_CLK), .Q(STATE[141]), .QN(n147) );
  DF3 STATE_reg_142_ ( .D(n604), .C(SYS_CLK), .Q(STATE[142]), .QN(n146) );
  DF3 STATE_reg_143_ ( .D(n603), .C(SYS_CLK), .Q(STATE[143]), .QN(n145) );
  DF3 STATE_reg_144_ ( .D(n602), .C(SYS_CLK), .Q(STATE[144]), .QN(n144) );
  DF3 STATE_reg_145_ ( .D(n601), .C(SYS_CLK), .Q(STATE[145]), .QN(n143) );
  DF3 STATE_reg_146_ ( .D(n600), .C(SYS_CLK), .Q(STATE[146]), .QN(n142) );
  DF3 STATE_reg_147_ ( .D(n599), .C(SYS_CLK), .Q(STATE[147]), .QN(n141) );
  DF3 STATE_reg_148_ ( .D(n598), .C(SYS_CLK), .Q(STATE[148]), .QN(n140) );
  DF3 STATE_reg_149_ ( .D(n597), .C(SYS_CLK), .Q(STATE[149]), .QN(n139) );
  DF3 STATE_reg_150_ ( .D(n596), .C(SYS_CLK), .Q(STATE[150]), .QN(n138) );
  DF3 STATE_reg_151_ ( .D(n595), .C(SYS_CLK), .Q(STATE[151]), .QN(n137) );
  DF3 STATE_reg_152_ ( .D(n594), .C(SYS_CLK), .Q(STATE[152]), .QN(n136) );
  DF3 STATE_reg_153_ ( .D(n593), .C(SYS_CLK), .Q(STATE[153]), .QN(n135) );
  DF3 STATE_reg_154_ ( .D(n592), .C(SYS_CLK), .Q(STATE[154]), .QN(n134) );
  DF3 STATE_reg_155_ ( .D(n591), .C(SYS_CLK), .Q(STATE[155]), .QN(n133) );
  DF3 STATE_reg_156_ ( .D(n590), .C(SYS_CLK), .Q(STATE[156]), .QN(n132) );
  DF3 STATE_reg_157_ ( .D(n589), .C(SYS_CLK), .Q(STATE[157]), .QN(n131) );
  DF3 STATE_reg_158_ ( .D(n588), .C(SYS_CLK), .Q(STATE[158]), .QN(n130) );
  DF3 STATE_reg_159_ ( .D(n587), .C(SYS_CLK), .Q(STATE[159]), .QN(n129) );
  DF3 STATE_reg_160_ ( .D(n586), .C(SYS_CLK), .Q(STATE[160]), .QN(n128) );
  DF3 STATE_reg_161_ ( .D(n585), .C(SYS_CLK), .Q(STATE[161]), .QN(n127) );
  DF3 STATE_reg_162_ ( .D(n584), .C(SYS_CLK), .Q(STATE[162]), .QN(n126) );
  DF3 STATE_reg_163_ ( .D(n583), .C(SYS_CLK), .Q(STATE[163]), .QN(n125) );
  DF3 STATE_reg_164_ ( .D(n582), .C(SYS_CLK), .Q(STATE[164]), .QN(n124) );
  DF3 STATE_reg_165_ ( .D(n581), .C(SYS_CLK), .Q(STATE[165]), .QN(n123) );
  DF3 STATE_reg_166_ ( .D(n580), .C(SYS_CLK), .Q(STATE[166]), .QN(n122) );
  DF3 STATE_reg_167_ ( .D(n579), .C(SYS_CLK), .Q(STATE[167]), .QN(n121) );
  DF3 STATE_reg_168_ ( .D(n578), .C(SYS_CLK), .Q(STATE[168]), .QN(n120) );
  DF3 STATE_reg_169_ ( .D(n577), .C(SYS_CLK), .Q(STATE[169]), .QN(n119) );
  DF3 STATE_reg_170_ ( .D(n576), .C(SYS_CLK), .Q(STATE[170]), .QN(n118) );
  DF3 STATE_reg_171_ ( .D(n575), .C(SYS_CLK), .Q(STATE[171]), .QN(n117) );
  DF3 STATE_reg_172_ ( .D(n574), .C(SYS_CLK), .QN(n116) );
  DF3 STATE_reg_173_ ( .D(n573), .C(SYS_CLK), .QN(n115) );
  DF3 STATE_reg_174_ ( .D(n572), .C(SYS_CLK), .QN(n114) );
  DF3 STATE_reg_175_ ( .D(n571), .C(SYS_CLK), .Q(STATE[175]), .QN(n113) );
  DF3 STATE_reg_176_ ( .D(n785), .C(SYS_CLK), .Q(STATE[176]) );
  DF3 STATE_reg_177_ ( .D(n784), .C(SYS_CLK), .Q(STATE[177]) );
  DF3 STATE_reg_178_ ( .D(n786), .C(SYS_CLK), .Q(STATE[178]) );
  DF3 STATE_reg_179_ ( .D(n787), .C(SYS_CLK), .Q(STATE[179]), .QN(n109) );
  DF3 STATE_reg_180_ ( .D(n570), .C(SYS_CLK), .QN(n108) );
  DF3 STATE_reg_181_ ( .D(n569), .C(SYS_CLK), .QN(n107) );
  DF3 STATE_reg_182_ ( .D(n568), .C(SYS_CLK), .QN(n106) );
  DF3 STATE_reg_183_ ( .D(n567), .C(SYS_CLK), .QN(n105) );
  DF3 STATE_reg_184_ ( .D(n566), .C(SYS_CLK), .QN(n104) );
  DF3 STATE_reg_185_ ( .D(n565), .C(SYS_CLK), .QN(n103) );
  DF3 STATE_reg_186_ ( .D(n564), .C(SYS_CLK), .QN(n102) );
  DF3 STATE_reg_187_ ( .D(n563), .C(SYS_CLK), .QN(n101) );
  DF3 STATE_reg_188_ ( .D(n562), .C(SYS_CLK), .QN(n100) );
  DF3 STATE_reg_189_ ( .D(n561), .C(SYS_CLK), .QN(n99) );
  DF3 STATE_reg_190_ ( .D(n560), .C(SYS_CLK), .QN(n98) );
  DF3 STATE_reg_191_ ( .D(n559), .C(SYS_CLK), .QN(n97) );
  DF3 STATE_reg_192_ ( .D(n558), .C(SYS_CLK), .QN(n96) );
  DF3 STATE_reg_193_ ( .D(n557), .C(SYS_CLK), .QN(n95) );
  DF3 STATE_reg_194_ ( .D(n556), .C(SYS_CLK), .QN(n94) );
  DF3 STATE_reg_195_ ( .D(n555), .C(SYS_CLK), .QN(n93) );
  DF3 STATE_reg_196_ ( .D(n554), .C(SYS_CLK), .QN(n92) );
  DF3 STATE_reg_197_ ( .D(n553), .C(SYS_CLK), .QN(n91) );
  DF3 STATE_reg_198_ ( .D(n552), .C(SYS_CLK), .QN(n90) );
  DF3 STATE_reg_199_ ( .D(n551), .C(SYS_CLK), .QN(n89) );
  DF3 STATE_reg_200_ ( .D(n550), .C(SYS_CLK), .QN(n88) );
  DF3 STATE_reg_201_ ( .D(n549), .C(SYS_CLK), .QN(n87) );
  DF3 STATE_reg_202_ ( .D(n548), .C(SYS_CLK), .QN(n86) );
  DF3 STATE_reg_203_ ( .D(n547), .C(SYS_CLK), .QN(n85) );
  DF3 STATE_reg_204_ ( .D(n546), .C(SYS_CLK), .QN(n84) );
  DF3 STATE_reg_205_ ( .D(n545), .C(SYS_CLK), .QN(n83) );
  DF3 STATE_reg_206_ ( .D(n544), .C(SYS_CLK), .QN(n82) );
  DF3 STATE_reg_207_ ( .D(n543), .C(SYS_CLK), .QN(n81) );
  DF3 STATE_reg_208_ ( .D(n542), .C(SYS_CLK), .QN(n80) );
  DF3 STATE_reg_209_ ( .D(n541), .C(SYS_CLK), .QN(n79) );
  DF3 STATE_reg_210_ ( .D(n540), .C(SYS_CLK), .QN(n78) );
  DF3 STATE_reg_211_ ( .D(n539), .C(SYS_CLK), .QN(n77) );
  DF3 STATE_reg_212_ ( .D(n538), .C(SYS_CLK), .QN(n76) );
  DF3 STATE_reg_213_ ( .D(n537), .C(SYS_CLK), .QN(n75) );
  DF3 STATE_reg_214_ ( .D(n536), .C(SYS_CLK), .QN(n74) );
  DF3 STATE_reg_215_ ( .D(n535), .C(SYS_CLK), .QN(n73) );
  DF3 STATE_reg_216_ ( .D(n534), .C(SYS_CLK), .QN(n72) );
  DF3 STATE_reg_217_ ( .D(n533), .C(SYS_CLK), .QN(n71) );
  DF3 STATE_reg_218_ ( .D(n532), .C(SYS_CLK), .QN(n70) );
  DF3 STATE_reg_219_ ( .D(n531), .C(SYS_CLK), .QN(n69) );
  DF3 STATE_reg_220_ ( .D(n530), .C(SYS_CLK), .QN(n68) );
  DF3 STATE_reg_221_ ( .D(n529), .C(SYS_CLK), .QN(n67) );
  DF3 STATE_reg_222_ ( .D(n528), .C(SYS_CLK), .QN(n66) );
  DF3 STATE_reg_223_ ( .D(n527), .C(SYS_CLK), .QN(n65) );
  DF3 STATE_reg_224_ ( .D(n526), .C(SYS_CLK), .QN(n64) );
  DF3 STATE_reg_225_ ( .D(n525), .C(SYS_CLK), .QN(n63) );
  DF3 STATE_reg_226_ ( .D(n524), .C(SYS_CLK), .QN(n62) );
  DF3 STATE_reg_227_ ( .D(n523), .C(SYS_CLK), .QN(n61) );
  DF3 STATE_reg_228_ ( .D(n522), .C(SYS_CLK), .QN(n60) );
  DF3 STATE_reg_229_ ( .D(n521), .C(SYS_CLK), .QN(n59) );
  DF3 STATE_reg_230_ ( .D(n520), .C(SYS_CLK), .QN(n58) );
  DF3 STATE_reg_231_ ( .D(n519), .C(SYS_CLK), .QN(n57) );
  DF3 STATE_reg_232_ ( .D(n518), .C(SYS_CLK), .QN(n56) );
  DF3 STATE_reg_233_ ( .D(n517), .C(SYS_CLK), .QN(n55) );
  DF3 STATE_reg_234_ ( .D(n516), .C(SYS_CLK), .QN(n54) );
  DF3 STATE_reg_235_ ( .D(n515), .C(SYS_CLK), .QN(n53) );
  DF3 STATE_reg_236_ ( .D(n514), .C(SYS_CLK), .QN(n52) );
  DF3 STATE_reg_237_ ( .D(n513), .C(SYS_CLK), .QN(n51) );
  DF3 STATE_reg_238_ ( .D(n512), .C(SYS_CLK), .QN(n50) );
  DF3 STATE_reg_239_ ( .D(n511), .C(SYS_CLK), .QN(n49) );
  DF3 STATE_reg_240_ ( .D(n510), .C(SYS_CLK), .QN(n48) );
  DF3 STATE_reg_241_ ( .D(n509), .C(SYS_CLK), .QN(n47) );
  DF3 STATE_reg_242_ ( .D(n508), .C(SYS_CLK), .Q(STATE[242]), .QN(n46) );
  DF3 STATE_reg_243_ ( .D(n507), .C(SYS_CLK), .QN(n45) );
  DF3 STATE_reg_244_ ( .D(n506), .C(SYS_CLK), .QN(n44) );
  DF3 STATE_reg_245_ ( .D(n505), .C(SYS_CLK), .QN(n43) );
  DF3 STATE_reg_246_ ( .D(n504), .C(SYS_CLK), .QN(n42) );
  DF3 STATE_reg_247_ ( .D(n503), .C(SYS_CLK), .QN(n41) );
  DF3 STATE_reg_248_ ( .D(n502), .C(SYS_CLK), .QN(n40) );
  DF3 STATE_reg_249_ ( .D(n501), .C(SYS_CLK), .QN(n39) );
  DF3 STATE_reg_250_ ( .D(n500), .C(SYS_CLK), .QN(n38) );
  DF3 STATE_reg_251_ ( .D(n499), .C(SYS_CLK), .QN(n37) );
  DF3 STATE_reg_252_ ( .D(n498), .C(SYS_CLK), .QN(n36) );
  DF3 STATE_reg_253_ ( .D(n497), .C(SYS_CLK), .QN(n35) );
  DF3 STATE_reg_254_ ( .D(n496), .C(SYS_CLK), .QN(n34) );
  DF3 STATE_reg_255_ ( .D(n495), .C(SYS_CLK), .QN(n33) );
  DF3 STATE_reg_256_ ( .D(n494), .C(SYS_CLK), .QN(n32) );
  DF3 STATE_reg_257_ ( .D(n493), .C(SYS_CLK), .QN(n31) );
  DF3 STATE_reg_258_ ( .D(n492), .C(SYS_CLK), .QN(n30) );
  DF3 STATE_reg_259_ ( .D(n491), .C(SYS_CLK), .QN(n29) );
  DF3 STATE_reg_260_ ( .D(n490), .C(SYS_CLK), .QN(n28) );
  DF3 STATE_reg_261_ ( .D(n489), .C(SYS_CLK), .QN(n27) );
  DF3 STATE_reg_262_ ( .D(n488), .C(SYS_CLK), .QN(n26) );
  DF3 STATE_reg_263_ ( .D(n487), .C(SYS_CLK), .Q(STATE[263]), .QN(n24) );
  DF3 STATE_reg_264_ ( .D(n486), .C(SYS_CLK), .QN(n23) );
  DF3 STATE_reg_265_ ( .D(n485), .C(SYS_CLK), .QN(n22) );
  DF3 STATE_reg_266_ ( .D(n484), .C(SYS_CLK), .QN(n21) );
  DF3 STATE_reg_267_ ( .D(n483), .C(SYS_CLK), .QN(n20) );
  DF3 STATE_reg_268_ ( .D(n482), .C(SYS_CLK), .QN(n19) );
  DF3 STATE_reg_269_ ( .D(n481), .C(SYS_CLK), .QN(n18) );
  DF3 STATE_reg_270_ ( .D(n480), .C(SYS_CLK), .QN(n17) );
  DF3 STATE_reg_271_ ( .D(n479), .C(SYS_CLK), .QN(n16) );
  DF3 STATE_reg_272_ ( .D(n478), .C(SYS_CLK), .QN(n15) );
  DF3 STATE_reg_273_ ( .D(n477), .C(SYS_CLK), .QN(n14) );
  DF3 STATE_reg_274_ ( .D(n476), .C(SYS_CLK), .QN(n13) );
  DF3 STATE_reg_275_ ( .D(n475), .C(SYS_CLK), .QN(n12) );
  DF3 STATE_reg_276_ ( .D(n474), .C(SYS_CLK), .QN(n11) );
  DF3 STATE_reg_277_ ( .D(n473), .C(SYS_CLK), .QN(n10) );
  DF3 STATE_reg_278_ ( .D(n472), .C(SYS_CLK), .QN(n9) );
  DF3 STATE_reg_279_ ( .D(n471), .C(SYS_CLK), .QN(n8) );
  DF3 STATE_reg_280_ ( .D(n470), .C(SYS_CLK), .QN(n7) );
  DF3 STATE_reg_281_ ( .D(n469), .C(SYS_CLK), .QN(n6) );
  DF3 STATE_reg_282_ ( .D(n468), .C(SYS_CLK), .QN(n5) );
  DF3 STATE_reg_283_ ( .D(n467), .C(SYS_CLK), .QN(n4) );
  DF3 STATE_reg_284_ ( .D(n466), .C(SYS_CLK), .QN(n3) );
  DF3 STATE_reg_285_ ( .D(n465), .C(SYS_CLK), .Q(STATE[285]), .QN(n2) );
  DF3 STATE_reg_286_ ( .D(n464), .C(SYS_CLK), .Q(STATE[286]), .QN(n1) );
  DF3 STATE_reg_287_ ( .D(n463), .C(SYS_CLK), .Q(STATE[287]) );
  XOR21 U474 ( .A(STATE[68]), .B(N305), .Q(n750) );
  XOR21 U477 ( .A(STATE[65]), .B(N301), .Q(n748) );
  XOR21 U480 ( .A(STATE[161]), .B(N303), .Q(n746) );
  XOR21 U479 ( .A(STATE[263]), .B(STATE[176]), .Q(n747) );
  XOR21 U481 ( .A(n747), .B(n746), .Q(t2) );
  XOR21 U468 ( .A(STATE[287]), .B(STATE[242]), .Q(n755) );
  XOR21 U469 ( .A(STATE[176]), .B(STATE[161]), .Q(n754) );
  XOR21 U471 ( .A(n755), .B(n754), .Q(n752) );
  XOR21 U470 ( .A(STATE[92]), .B(STATE[65]), .Q(n753) );
  XOR21 U472 ( .A(n753), .B(n752), .Q(KEY_OUT) );
  NOR20 U4 ( .A(n289), .B(n782), .Q(n298) );
  INV2 U6 ( .A(n111), .Q(n112) );
  NOR20 U8 ( .A(n788), .B(CNTRL[0]), .Q(n294) );
  CLKBU2 U114 ( .A(n112), .Q(n782) );
  AOI221 U115 ( .A(IV[7]), .B(n779), .C(t1), .D(n767), .Q(n381) );
  AOI221 U116 ( .A(KEY[7]), .B(n779), .C(t3), .D(n768), .Q(n462) );
  INV3 U117 ( .A(n777), .Q(n765) );
  INV3 U122 ( .A(n777), .Q(n766) );
  INV3 U124 ( .A(n776), .Q(n767) );
  INV3 U126 ( .A(n290), .Q(n768) );
  BUF2 U128 ( .A(n776), .Q(n775) );
  BUF2 U130 ( .A(n777), .Q(n774) );
  BUF2 U132 ( .A(n776), .Q(n773) );
  BUF2 U134 ( .A(n777), .Q(n772) );
  BUF2 U136 ( .A(n777), .Q(n771) );
  BUF2 U138 ( .A(n776), .Q(n770) );
  BUF2 U140 ( .A(n777), .Q(n769) );
  BUF2 U142 ( .A(n756), .Q(n759) );
  BUF2 U144 ( .A(n751), .Q(n761) );
  BUF2 U146 ( .A(n749), .Q(n760) );
  BUF2 U148 ( .A(n751), .Q(n762) );
  BUF2 U150 ( .A(n758), .Q(n763) );
  BUF2 U152 ( .A(n758), .Q(n764) );
  INV3 U154 ( .A(n291), .Q(n776) );
  INV3 U156 ( .A(n291), .Q(n777) );
  INV3 U158 ( .A(n290), .Q(n291) );
  BUF2 U160 ( .A(n196), .Q(n758) );
  BUF2 U162 ( .A(n196), .Q(n757) );
  BUF2 U164 ( .A(n196), .Q(n756) );
  BUF2 U166 ( .A(n196), .Q(n749) );
  BUF2 U168 ( .A(n196), .Q(n751) );
  INV3 U170 ( .A(n298), .Q(n290) );
  BUF2 U172 ( .A(n112), .Q(n781) );
  BUF2 U174 ( .A(n781), .Q(n780) );
  BUF2 U176 ( .A(n778), .Q(n779) );
  BUF2 U178 ( .A(n112), .Q(n778) );
  INV3 U180 ( .A(n196), .Q(n289) );
  AOI221 U182 ( .A(KEY[3]), .B(n112), .C(STATE[3]), .D(n768), .Q(n458) );
  AOI221 U184 ( .A(KEY[4]), .B(n112), .C(STATE[2]), .D(n768), .Q(n459) );
  AOI221 U186 ( .A(KEY[5]), .B(n112), .C(STATE[1]), .D(n768), .Q(n460) );
  AOI221 U188 ( .A(KEY[6]), .B(n112), .C(STATE[0]), .D(n768), .Q(n461) );
  XNR21 U190 ( .A(n25), .B(n750), .Q(t3) );
  XNR21 U192 ( .A(STATE[287]), .B(STATE[242]), .Q(n25) );
  AOI221 U194 ( .A(IV[72]), .B(n778), .C(STATE[171]), .D(n768), .Q(n302) );
  AOI221 U196 ( .A(KEY[72]), .B(n778), .C(STATE[78]), .D(n767), .Q(n383) );
  AOI221 U198 ( .A(IV[73]), .B(n782), .C(STATE[170]), .D(n768), .Q(n303) );
  AOI221 U200 ( .A(IV[74]), .B(n781), .C(STATE[169]), .D(n768), .Q(n304) );
  AOI221 U202 ( .A(IV[75]), .B(n778), .C(STATE[168]), .D(n765), .Q(n305) );
  AOI221 U204 ( .A(IV[76]), .B(n782), .C(STATE[167]), .D(n768), .Q(n306) );
  AOI221 U206 ( .A(IV[77]), .B(n782), .C(STATE[166]), .D(n768), .Q(n307) );
  AOI221 U208 ( .A(IV[78]), .B(n781), .C(STATE[165]), .D(n298), .Q(n308) );
  AOI221 U210 ( .A(IV[79]), .B(n778), .C(STATE[164]), .D(n767), .Q(n309) );
  AOI221 U212 ( .A(IV[64]), .B(n781), .C(STATE[163]), .D(n767), .Q(n310) );
  AOI221 U214 ( .A(IV[65]), .B(n782), .C(STATE[162]), .D(n768), .Q(n311) );
  AOI221 U216 ( .A(IV[66]), .B(n782), .C(STATE[161]), .D(n768), .Q(n312) );
  AOI221 U218 ( .A(IV[67]), .B(n782), .C(STATE[160]), .D(n768), .Q(n313) );
  AOI221 U220 ( .A(IV[68]), .B(n782), .C(STATE[159]), .D(n765), .Q(n314) );
  AOI221 U222 ( .A(IV[69]), .B(n782), .C(STATE[158]), .D(n765), .Q(n315) );
  AOI221 U224 ( .A(IV[70]), .B(n782), .C(STATE[157]), .D(n765), .Q(n316) );
  AOI221 U226 ( .A(IV[71]), .B(n782), .C(STATE[156]), .D(n765), .Q(n317) );
  AOI221 U228 ( .A(IV[56]), .B(n782), .C(STATE[155]), .D(n765), .Q(n318) );
  AOI221 U230 ( .A(IV[57]), .B(n782), .C(STATE[154]), .D(n765), .Q(n319) );
  AOI221 U232 ( .A(IV[58]), .B(n782), .C(STATE[153]), .D(n765), .Q(n320) );
  AOI221 U234 ( .A(IV[59]), .B(n782), .C(STATE[152]), .D(n765), .Q(n321) );
  AOI221 U236 ( .A(IV[60]), .B(n782), .C(STATE[151]), .D(n765), .Q(n322) );
  AOI221 U238 ( .A(IV[61]), .B(n782), .C(STATE[150]), .D(n765), .Q(n323) );
  AOI221 U240 ( .A(IV[62]), .B(n782), .C(STATE[149]), .D(n765), .Q(n324) );
  AOI221 U242 ( .A(IV[63]), .B(n782), .C(STATE[148]), .D(n765), .Q(n325) );
  AOI221 U244 ( .A(IV[48]), .B(n782), .C(STATE[147]), .D(n765), .Q(n326) );
  AOI221 U246 ( .A(IV[49]), .B(n782), .C(STATE[146]), .D(n766), .Q(n327) );
  AOI221 U248 ( .A(IV[50]), .B(n782), .C(STATE[145]), .D(n766), .Q(n328) );
  AOI221 U250 ( .A(IV[51]), .B(n779), .C(STATE[144]), .D(n766), .Q(n329) );
  AOI221 U252 ( .A(IV[52]), .B(n780), .C(STATE[143]), .D(n766), .Q(n330) );
  AOI221 U254 ( .A(IV[53]), .B(n779), .C(STATE[142]), .D(n766), .Q(n331) );
  AOI221 U256 ( .A(IV[54]), .B(n780), .C(STATE[141]), .D(n766), .Q(n332) );
  AOI221 U258 ( .A(IV[55]), .B(n779), .C(STATE[140]), .D(n766), .Q(n333) );
  AOI221 U260 ( .A(IV[40]), .B(n780), .C(STATE[139]), .D(n766), .Q(n334) );
  AOI221 U262 ( .A(IV[41]), .B(n779), .C(STATE[138]), .D(n766), .Q(n335) );
  AOI221 U264 ( .A(IV[42]), .B(n780), .C(STATE[137]), .D(n766), .Q(n336) );
  AOI221 U266 ( .A(IV[43]), .B(n779), .C(STATE[136]), .D(n766), .Q(n337) );
  AOI221 U268 ( .A(IV[44]), .B(n780), .C(STATE[135]), .D(n767), .Q(n338) );
  AOI221 U270 ( .A(IV[45]), .B(n112), .C(STATE[134]), .D(n766), .Q(n339) );
  AOI221 U272 ( .A(IV[46]), .B(n112), .C(STATE[133]), .D(n766), .Q(n340) );
  AOI221 U274 ( .A(IV[47]), .B(n294), .C(STATE[132]), .D(n765), .Q(n341) );
  AOI221 U276 ( .A(IV[32]), .B(n294), .C(STATE[131]), .D(n766), .Q(n342) );
  AOI221 U278 ( .A(IV[33]), .B(n294), .C(STATE[130]), .D(n765), .Q(n343) );
  AOI221 U280 ( .A(IV[34]), .B(n294), .C(STATE[129]), .D(n766), .Q(n344) );
  AOI221 U281 ( .A(IV[35]), .B(n294), .C(STATE[128]), .D(n765), .Q(n345) );
  AOI221 U295 ( .A(IV[36]), .B(n781), .C(STATE[127]), .D(n766), .Q(n346) );
  AOI221 U297 ( .A(IV[37]), .B(n781), .C(STATE[126]), .D(n765), .Q(n347) );
  AOI221 U299 ( .A(IV[38]), .B(n781), .C(STATE[125]), .D(n766), .Q(n348) );
  AOI221 U301 ( .A(IV[39]), .B(n781), .C(STATE[124]), .D(n765), .Q(n349) );
  AOI221 U303 ( .A(IV[24]), .B(n781), .C(STATE[123]), .D(n766), .Q(n350) );
  AOI221 U305 ( .A(IV[25]), .B(n781), .C(STATE[122]), .D(n765), .Q(n351) );
  AOI221 U307 ( .A(IV[26]), .B(n781), .C(STATE[121]), .D(n766), .Q(n352) );
  AOI221 U309 ( .A(IV[27]), .B(n781), .C(STATE[120]), .D(n765), .Q(n353) );
  AOI221 U311 ( .A(IV[28]), .B(n781), .C(STATE[119]), .D(n298), .Q(n354) );
  AOI221 U313 ( .A(IV[29]), .B(n781), .C(STATE[118]), .D(n298), .Q(n355) );
  AOI221 U315 ( .A(IV[30]), .B(n781), .C(STATE[117]), .D(n291), .Q(n356) );
  AOI221 U317 ( .A(IV[31]), .B(n781), .C(STATE[116]), .D(n291), .Q(n357) );
  AOI221 U319 ( .A(IV[16]), .B(n781), .C(STATE[115]), .D(n291), .Q(n358) );
  AOI221 U321 ( .A(IV[17]), .B(n781), .C(STATE[114]), .D(n291), .Q(n359) );
  AOI221 U323 ( .A(IV[18]), .B(n781), .C(STATE[113]), .D(n291), .Q(n360) );
  AOI221 U325 ( .A(IV[19]), .B(n781), .C(STATE[112]), .D(n291), .Q(n361) );
  AOI221 U327 ( .A(IV[20]), .B(n781), .C(STATE[111]), .D(n291), .Q(n362) );
  AOI221 U329 ( .A(IV[21]), .B(n780), .C(STATE[110]), .D(n765), .Q(n363) );
  AOI221 U331 ( .A(IV[22]), .B(n780), .C(STATE[109]), .D(n291), .Q(n364) );
  AOI221 U333 ( .A(IV[23]), .B(n780), .C(STATE[108]), .D(n291), .Q(n365) );
  AOI221 U335 ( .A(IV[8]), .B(n780), .C(STATE[107]), .D(n291), .Q(n366) );
  AOI221 U337 ( .A(IV[9]), .B(n780), .C(STATE[106]), .D(n768), .Q(n367) );
  AOI221 U339 ( .A(IV[10]), .B(n780), .C(STATE[105]), .D(n768), .Q(n368) );
  AOI221 U341 ( .A(IV[11]), .B(n780), .C(STATE[104]), .D(n768), .Q(n369) );
  AOI221 U343 ( .A(IV[12]), .B(n780), .C(STATE[103]), .D(n768), .Q(n370) );
  AOI221 U345 ( .A(IV[13]), .B(n780), .C(STATE[102]), .D(n768), .Q(n371) );
  AOI221 U347 ( .A(IV[14]), .B(n780), .C(STATE[101]), .D(n768), .Q(n372) );
  AOI221 U349 ( .A(IV[15]), .B(n780), .C(STATE[100]), .D(n768), .Q(n373) );
  AOI221 U351 ( .A(IV[0]), .B(n780), .C(STATE[99]), .D(n768), .Q(n374) );
  AOI221 U353 ( .A(IV[1]), .B(n780), .C(STATE[98]), .D(n291), .Q(n375) );
  AOI221 U355 ( .A(IV[2]), .B(n780), .C(STATE[97]), .D(n767), .Q(n376) );
  AOI221 U357 ( .A(IV[3]), .B(n780), .C(STATE[96]), .D(n765), .Q(n377) );
  AOI221 U359 ( .A(IV[4]), .B(n780), .C(STATE[95]), .D(n766), .Q(n378) );
  AOI221 U361 ( .A(IV[5]), .B(n780), .C(STATE[94]), .D(n291), .Q(n379) );
  AOI221 U363 ( .A(IV[6]), .B(n782), .C(STATE[93]), .D(n767), .Q(n380) );
  XNR21 U365 ( .A(n110), .B(n748), .Q(t1) );
  XNR21 U367 ( .A(STATE[170]), .B(STATE[92]), .Q(n110) );
  AOI221 U369 ( .A(KEY[76]), .B(n781), .C(STATE[74]), .D(n767), .Q(n387) );
  AOI221 U371 ( .A(KEY[77]), .B(n780), .C(STATE[73]), .D(n767), .Q(n388) );
  AOI221 U373 ( .A(KEY[78]), .B(n779), .C(STATE[72]), .D(n767), .Q(n389) );
  AOI221 U375 ( .A(KEY[79]), .B(n782), .C(STATE[71]), .D(n767), .Q(n390) );
  AOI221 U377 ( .A(KEY[64]), .B(n780), .C(STATE[70]), .D(n767), .Q(n391) );
  AOI221 U379 ( .A(KEY[65]), .B(n779), .C(STATE[69]), .D(n767), .Q(n392) );
  AOI221 U381 ( .A(KEY[66]), .B(n780), .C(STATE[68]), .D(n768), .Q(n393) );
  AOI221 U383 ( .A(KEY[67]), .B(n780), .C(STATE[67]), .D(n767), .Q(n394) );
  AOI221 U385 ( .A(KEY[68]), .B(n779), .C(STATE[66]), .D(n768), .Q(n395) );
  AOI221 U387 ( .A(KEY[69]), .B(n779), .C(STATE[65]), .D(n766), .Q(n396) );
  AOI221 U389 ( .A(KEY[70]), .B(n780), .C(STATE[64]), .D(n765), .Q(n397) );
  AOI221 U391 ( .A(KEY[71]), .B(n779), .C(STATE[63]), .D(n766), .Q(n398) );
  AOI221 U393 ( .A(KEY[56]), .B(n779), .C(STATE[62]), .D(n767), .Q(n399) );
  AOI221 U395 ( .A(KEY[57]), .B(n779), .C(STATE[61]), .D(n291), .Q(n400) );
  AOI221 U397 ( .A(KEY[58]), .B(n779), .C(STATE[60]), .D(n768), .Q(n401) );
  AOI221 U399 ( .A(KEY[59]), .B(n779), .C(STATE[59]), .D(n291), .Q(n402) );
  AOI221 U401 ( .A(KEY[60]), .B(n779), .C(STATE[58]), .D(n768), .Q(n403) );
  AOI221 U403 ( .A(KEY[61]), .B(n779), .C(STATE[57]), .D(n765), .Q(n404) );
  AOI221 U405 ( .A(KEY[62]), .B(n779), .C(STATE[56]), .D(n291), .Q(n405) );
  AOI221 U407 ( .A(KEY[63]), .B(n779), .C(STATE[55]), .D(n767), .Q(n406) );
  AOI221 U409 ( .A(KEY[48]), .B(n779), .C(STATE[54]), .D(n291), .Q(n407) );
  AOI221 U411 ( .A(KEY[49]), .B(n779), .C(STATE[53]), .D(n765), .Q(n408) );
  AOI221 U413 ( .A(KEY[50]), .B(n779), .C(STATE[52]), .D(n766), .Q(n409) );
  AOI221 U415 ( .A(KEY[51]), .B(n779), .C(STATE[51]), .D(n767), .Q(n410) );
  AOI221 U417 ( .A(KEY[52]), .B(n779), .C(STATE[50]), .D(n767), .Q(n411) );
  AOI221 U419 ( .A(KEY[53]), .B(n779), .C(STATE[49]), .D(n768), .Q(n412) );
  AOI221 U421 ( .A(KEY[54]), .B(n779), .C(STATE[48]), .D(n766), .Q(n413) );
  AOI221 U423 ( .A(KEY[55]), .B(n779), .C(STATE[47]), .D(n768), .Q(n414) );
  AOI221 U425 ( .A(KEY[40]), .B(n778), .C(STATE[46]), .D(n767), .Q(n415) );
  AOI221 U427 ( .A(KEY[41]), .B(n778), .C(STATE[45]), .D(n765), .Q(n416) );
  AOI221 U429 ( .A(KEY[42]), .B(n778), .C(STATE[44]), .D(n766), .Q(n417) );
  AOI221 U431 ( .A(KEY[43]), .B(n778), .C(STATE[43]), .D(n291), .Q(n418) );
  AOI221 U433 ( .A(KEY[44]), .B(n778), .C(STATE[42]), .D(n765), .Q(n419) );
  AOI221 U435 ( .A(KEY[45]), .B(n778), .C(STATE[41]), .D(n291), .Q(n420) );
  AOI221 U437 ( .A(KEY[46]), .B(n778), .C(STATE[40]), .D(n768), .Q(n421) );
  AOI221 U439 ( .A(KEY[47]), .B(n778), .C(STATE[39]), .D(n766), .Q(n422) );
  AOI221 U441 ( .A(KEY[32]), .B(n778), .C(STATE[38]), .D(n291), .Q(n423) );
  AOI221 U443 ( .A(KEY[33]), .B(n778), .C(STATE[37]), .D(n291), .Q(n424) );
  AOI221 U445 ( .A(KEY[34]), .B(n778), .C(STATE[36]), .D(n768), .Q(n425) );
  AOI221 U447 ( .A(KEY[35]), .B(n778), .C(STATE[35]), .D(n298), .Q(n426) );
  AOI221 U449 ( .A(KEY[36]), .B(n778), .C(STATE[34]), .D(n291), .Q(n427) );
  AOI221 U451 ( .A(KEY[37]), .B(n778), .C(STATE[33]), .D(n766), .Q(n428) );
  AOI221 U453 ( .A(KEY[38]), .B(n778), .C(STATE[32]), .D(n298), .Q(n429) );
  AOI221 U454 ( .A(KEY[39]), .B(n778), .C(STATE[31]), .D(n766), .Q(n430) );
  AOI221 U455 ( .A(KEY[24]), .B(n778), .C(STATE[30]), .D(n768), .Q(n431) );
  AOI221 U456 ( .A(KEY[25]), .B(n778), .C(STATE[29]), .D(n767), .Q(n432) );
  AOI221 U457 ( .A(KEY[26]), .B(n782), .C(STATE[28]), .D(n768), .Q(n433) );
  AOI221 U458 ( .A(KEY[27]), .B(n778), .C(STATE[27]), .D(n768), .Q(n434) );
  AOI221 U459 ( .A(KEY[28]), .B(n782), .C(STATE[26]), .D(n768), .Q(n435) );
  AOI221 U460 ( .A(KEY[29]), .B(n781), .C(STATE[25]), .D(n765), .Q(n436) );
  AOI221 U461 ( .A(KEY[30]), .B(n778), .C(STATE[24]), .D(n298), .Q(n437) );
  AOI221 U462 ( .A(KEY[31]), .B(n782), .C(STATE[23]), .D(n768), .Q(n438) );
  AOI221 U463 ( .A(KEY[16]), .B(n781), .C(STATE[22]), .D(n765), .Q(n439) );
  AOI221 U464 ( .A(KEY[17]), .B(n781), .C(STATE[21]), .D(n767), .Q(n440) );
  AOI221 U465 ( .A(KEY[18]), .B(n778), .C(STATE[20]), .D(n765), .Q(n441) );
  AOI221 U466 ( .A(KEY[19]), .B(n781), .C(STATE[19]), .D(n766), .Q(n442) );
  AOI221 U467 ( .A(KEY[20]), .B(n778), .C(STATE[18]), .D(n291), .Q(n443) );
  AOI221 U473 ( .A(KEY[21]), .B(n782), .C(STATE[17]), .D(n768), .Q(n444) );
  AOI221 U475 ( .A(KEY[22]), .B(n781), .C(STATE[16]), .D(n768), .Q(n445) );
  AOI221 U476 ( .A(KEY[23]), .B(n778), .C(STATE[15]), .D(n768), .Q(n446) );
  AOI221 U478 ( .A(KEY[8]), .B(n782), .C(STATE[14]), .D(n768), .Q(n447) );
  AOI221 U482 ( .A(KEY[9]), .B(n781), .C(STATE[13]), .D(n768), .Q(n448) );
  AOI221 U483 ( .A(KEY[10]), .B(n112), .C(STATE[12]), .D(n768), .Q(n449) );
  AOI221 U484 ( .A(KEY[11]), .B(n112), .C(STATE[11]), .D(n768), .Q(n450) );
  AOI221 U485 ( .A(KEY[12]), .B(n112), .C(STATE[10]), .D(n768), .Q(n451) );
  AOI221 U486 ( .A(KEY[13]), .B(n112), .C(STATE[9]), .D(n766), .Q(n452) );
  AOI221 U487 ( .A(KEY[14]), .B(n112), .C(STATE[8]), .D(n291), .Q(n453) );
  AOI221 U488 ( .A(KEY[15]), .B(n112), .C(STATE[7]), .D(n766), .Q(n454) );
  AOI221 U489 ( .A(KEY[0]), .B(n112), .C(STATE[6]), .D(n767), .Q(n455) );
  AOI221 U490 ( .A(KEY[1]), .B(n112), .C(STATE[5]), .D(n765), .Q(n456) );
  AOI221 U491 ( .A(KEY[2]), .B(n112), .C(STATE[4]), .D(n766), .Q(n457) );
  AOI221 U492 ( .A(KEY[73]), .B(n779), .C(STATE[77]), .D(n767), .Q(n384) );
  AOI221 U493 ( .A(KEY[74]), .B(n780), .C(STATE[76]), .D(n767), .Q(n385) );
  AOI221 U494 ( .A(KEY[75]), .B(n780), .C(STATE[75]), .D(n767), .Q(n386) );
  INV3 U495 ( .A(n292), .Q(n196) );
  NOR21 U496 ( .A(CNTRL[0]), .B(n294), .Q(n292) );
  INV3 U497 ( .A(n294), .Q(n111) );
  INV3 U498 ( .A(CNTRL[1]), .Q(n788) );
  INV3 U499 ( .A(n301), .Q(n785) );
  AOI221 U500 ( .A(n289), .B(STATE[176]), .C(n768), .D(STATE[175]), .Q(n301)
         );
  INV3 U501 ( .A(n382), .Q(n783) );
  AOI221 U502 ( .A(n289), .B(STATE[92]), .C(n768), .D(STATE[91]), .Q(n382) );
  AOI211 U503 ( .A(STATE[287]), .B(n289), .C(n782), .Q(n293) );
  AOI211 U504 ( .A(STATE[286]), .B(n292), .C(n781), .Q(n295) );
  AOI211 U505 ( .A(STATE[285]), .B(n289), .C(n778), .Q(n296) );
  INV3 U506 ( .A(n297), .Q(n787) );
  AOI221 U507 ( .A(n289), .B(STATE[179]), .C(n768), .D(STATE[178]), .Q(n297)
         );
  INV3 U508 ( .A(n299), .Q(n786) );
  AOI221 U509 ( .A(n289), .B(STATE[178]), .C(n768), .D(STATE[177]), .Q(n299)
         );
  INV3 U510 ( .A(n300), .Q(n784) );
  AOI221 U511 ( .A(n289), .B(STATE[177]), .C(n768), .D(t2), .Q(n300) );
  NOR21 U512 ( .A(n113), .B(n114), .Q(N303) );
  NOR21 U513 ( .A(n197), .B(n198), .Q(N301) );
  NOR21 U514 ( .A(n1), .B(n2), .Q(N305) );
endmodule


module Trivium_Generator_vvect_DW01_inc_0 ( A, SUM );
  input [10:0] A;
  output [10:0] SUM;

  wire   [10:2] carry;

  ADD22 U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .S(SUM[9]) );
  ADD22 U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  ADD22 U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  ADD22 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  ADD22 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADD22 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADD22 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADD22 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADD22 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  INV3 U1 ( .A(A[0]), .Q(SUM[0]) );
  XOR20 U2 ( .A(carry[10]), .B(A[10]), .Q(SUM[10]) );
endmodule


module Trivium_Generator_vvect ( SYS_CLK, RST, PLAINTEXT_IN, CIPHERTEXT_OUT, 
        K_INPUT, IV_INPUT, PLNTXT_EN, CPHRTXT_RDY );
  input [79:0] K_INPUT;
  input [79:0] IV_INPUT;
  input SYS_CLK, RST, PLAINTEXT_IN, PLNTXT_EN;
  output CIPHERTEXT_OUT, CPHRTXT_RDY;
  wire   CORE_OUT, N21, N22, N23, N56, N57, N58, N59, N60, N61, N62, N63, N64,
         N65, N66, n15, n17, n18, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77;
  wire   [1:0] CORE_CNTRL;
  wire   [2:0] pr_state;
  wire   [10:0] INIT_COUNTER;

  OAI212 U32 ( .A(n50), .B(n23), .C(pr_state[0]), .Q(n49) );
  OAI212 U37 ( .A(n18), .B(n52), .C(n15), .Q(n51) );
  DF3 INIT_COUNTER_reg_0_ ( .D(n61), .C(SYS_CLK), .Q(INIT_COUNTER[0]) );
  DF3 pr_state_reg_0_ ( .D(N21), .C(SYS_CLK), .Q(pr_state[0]), .QN(n18) );
  DF3 pr_state_reg_1_ ( .D(N22), .C(SYS_CLK), .Q(pr_state[1]), .QN(n17) );
  DF3 pr_state_reg_2_ ( .D(N23), .C(SYS_CLK), .Q(pr_state[2]), .QN(n15) );
  DF3 INIT_COUNTER_reg_1_ ( .D(n71), .C(SYS_CLK), .Q(INIT_COUNTER[1]) );
  DF3 INIT_COUNTER_reg_2_ ( .D(n70), .C(SYS_CLK), .Q(INIT_COUNTER[2]) );
  DF3 INIT_COUNTER_reg_3_ ( .D(n69), .C(SYS_CLK), .Q(INIT_COUNTER[3]) );
  DF3 INIT_COUNTER_reg_4_ ( .D(n68), .C(SYS_CLK), .Q(INIT_COUNTER[4]) );
  DF3 INIT_COUNTER_reg_5_ ( .D(n67), .C(SYS_CLK), .Q(INIT_COUNTER[5]) );
  DF3 INIT_COUNTER_reg_6_ ( .D(n66), .C(SYS_CLK), .Q(INIT_COUNTER[6]) );
  DF3 INIT_COUNTER_reg_7_ ( .D(n65), .C(SYS_CLK), .Q(INIT_COUNTER[7]) );
  DF3 INIT_COUNTER_reg_8_ ( .D(n64), .C(SYS_CLK), .Q(INIT_COUNTER[8]) );
  DF3 INIT_COUNTER_reg_9_ ( .D(n63), .C(SYS_CLK), .Q(INIT_COUNTER[9]) );
  DF3 INIT_COUNTER_reg_10_ ( .D(n62), .C(SYS_CLK), .Q(INIT_COUNTER[10]) );
  DF3 CORE_CNTRL_reg_1_ ( .D(n73), .C(SYS_CLK), .Q(CORE_CNTRL[1]) );
  DF3 CORE_CNTRL_reg_0_ ( .D(n59), .C(SYS_CLK), .Q(CORE_CNTRL[0]) );
  DF3 CPHRTXT_RDY_reg ( .D(n58), .C(SYS_CLK), .Q(CPHRTXT_RDY) );
  DF3 CIPHERTEXT_OUT_reg ( .D(n57), .C(SYS_CLK), .Q(CIPHERTEXT_OUT) );
  TRIVIUM_CORE TRIV_CORE_GEN ( .SYS_CLK(SYS_CLK), .CNTRL(CORE_CNTRL), .KEY(
        K_INPUT), .IV(IV_INPUT), .KEY_OUT(CORE_OUT) );
  Trivium_Generator_vvect_DW01_inc_0 add_184 ( .A(INIT_COUNTER), .SUM({N66, 
        N65, N64, N63, N62, N61, N60, N59, N58, N57, N56}) );
  INV3 U62 ( .A(n32), .Q(n75) );
  NAND31 U63 ( .A(n33), .B(n34), .C(n35), .Q(n32) );
  NOR21 U64 ( .A(n35), .B(n23), .Q(n37) );
  NOR21 U65 ( .A(n23), .B(n29), .Q(n35) );
  INV3 U66 ( .A(n34), .Q(n76) );
  INV3 U67 ( .A(n33), .Q(n74) );
  INV3 U68 ( .A(n36), .Q(n62) );
  AOI221 U69 ( .A(n35), .B(INIT_COUNTER[10]), .C(n37), .D(N66), .Q(n36) );
  INV3 U70 ( .A(n38), .Q(n63) );
  AOI221 U71 ( .A(n35), .B(INIT_COUNTER[9]), .C(n37), .D(N65), .Q(n38) );
  INV3 U72 ( .A(n39), .Q(n64) );
  AOI221 U73 ( .A(n35), .B(INIT_COUNTER[8]), .C(n37), .D(N64), .Q(n39) );
  INV3 U74 ( .A(n40), .Q(n65) );
  AOI221 U75 ( .A(n35), .B(INIT_COUNTER[7]), .C(n37), .D(N63), .Q(n40) );
  INV3 U76 ( .A(n41), .Q(n66) );
  AOI221 U77 ( .A(n35), .B(INIT_COUNTER[6]), .C(n37), .D(N62), .Q(n41) );
  NOR21 U78 ( .A(pr_state[1]), .B(pr_state[2]), .Q(n23) );
  NOR31 U79 ( .A(n18), .B(pr_state[2]), .C(n17), .Q(n29) );
  INV3 U80 ( .A(n53), .Q(n72) );
  NAND41 U81 ( .A(INIT_COUNTER[0]), .B(INIT_COUNTER[1]), .C(n77), .D(n54), .Q(
        n53) );
  INV3 U82 ( .A(n56), .Q(n77) );
  NOR40 U83 ( .A(n55), .B(INIT_COUNTER[7]), .C(INIT_COUNTER[9]), .D(
        INIT_COUNTER[8]), .Q(n54) );
  OAI311 U84 ( .A(n30), .B(n23), .C(n74), .D(n31), .Q(n59) );
  NAND22 U85 ( .A(CORE_CNTRL[0]), .B(n75), .Q(n31) );
  OAI311 U86 ( .A(n18), .B(PLNTXT_EN), .C(n29), .D(n32), .Q(n30) );
  INV3 U87 ( .A(n28), .Q(n73) );
  AOI2111 U88 ( .A(n75), .B(CORE_CNTRL[1]), .C(n74), .D(n29), .Q(n28) );
  INV3 U89 ( .A(n47), .Q(n61) );
  AOI221 U90 ( .A(n35), .B(INIT_COUNTER[0]), .C(n37), .D(N56), .Q(n47) );
  NAND31 U91 ( .A(INIT_COUNTER[6]), .B(INIT_COUNTER[10]), .C(INIT_COUNTER[5]), 
        .Q(n55) );
  INV3 U92 ( .A(n44), .Q(n69) );
  AOI221 U93 ( .A(n35), .B(INIT_COUNTER[3]), .C(n37), .D(N59), .Q(n44) );
  INV3 U94 ( .A(n46), .Q(n71) );
  AOI221 U95 ( .A(n35), .B(INIT_COUNTER[1]), .C(n37), .D(N57), .Q(n46) );
  INV3 U96 ( .A(n45), .Q(n70) );
  AOI221 U97 ( .A(n35), .B(INIT_COUNTER[2]), .C(n37), .D(N58), .Q(n45) );
  AOI211 U98 ( .A(n34), .B(n51), .C(RST), .Q(N21) );
  NOR21 U99 ( .A(n72), .B(n17), .Q(n52) );
  OAI311 U100 ( .A(n22), .B(n23), .C(n24), .D(n25), .Q(n57) );
  NAND22 U101 ( .A(CIPHERTEXT_OUT), .B(n24), .Q(n25) );
  AOI311 U102 ( .A(PLNTXT_EN), .B(pr_state[0]), .C(n76), .D(n23), .Q(n24) );
  XNR21 U103 ( .A(PLAINTEXT_IN), .B(CORE_OUT), .Q(n22) );
  AOI211 U104 ( .A(n33), .B(n49), .C(RST), .Q(N22) );
  NOR21 U105 ( .A(pr_state[2]), .B(n72), .Q(n50) );
  INV3 U106 ( .A(n42), .Q(n67) );
  AOI221 U107 ( .A(n35), .B(INIT_COUNTER[5]), .C(n37), .D(N61), .Q(n42) );
  INV3 U108 ( .A(n43), .Q(n68) );
  AOI221 U109 ( .A(n35), .B(INIT_COUNTER[4]), .C(n37), .D(N60), .Q(n43) );
  NAND31 U110 ( .A(n18), .B(n15), .C(pr_state[1]), .Q(n33) );
  NAND31 U111 ( .A(INIT_COUNTER[2]), .B(INIT_COUNTER[4]), .C(INIT_COUNTER[3]), 
        .Q(n56) );
  NAND22 U112 ( .A(pr_state[2]), .B(n17), .Q(n34) );
  OAI311 U113 ( .A(n60), .B(n23), .C(n26), .D(n27), .Q(n58) );
  INV3 U114 ( .A(PLNTXT_EN), .Q(n60) );
  NAND22 U115 ( .A(CPHRTXT_RDY), .B(n26), .Q(n27) );
  AOI211 U116 ( .A(pr_state[0]), .B(n76), .C(n23), .Q(n26) );
  NOR21 U117 ( .A(RST), .B(n48), .Q(N23) );
  AOI211 U118 ( .A(n29), .B(n72), .C(n76), .Q(n48) );
endmodule

